module FPCategorical
#(parameter N = 8)
(
  input         clk,
  input         rst,
  input  [30:0] in_a,
  output [30:0] out_b
);


endmodule